// Lets say that the environment class was already there, and generator is
// a new component that needs to be included in the ENV.
class env;
  generator 	g0; 			      // Generate transactions
  driver 			d0; 			      // Driver to design
  monitor 		m0; 			      // Monitor from design
  scoreboard 	s0; 			      // Scoreboard connected to monitor
  mailbox 		scb_mbx; 		    // Top level mailbox for SCB <-> MON
  virtual bus_if 	m_bus_vif; 	// Virtual interface handle

  event drv_done;
  mailbox drv_mbx;

  function new();
    $display("T=%0t [Env] constructor", $time);
    d0 = new();
    m0 = new();
    s0 = new();
    scb_mbx = new();
    g0 = new();
    drv_mbx = new();
  endfunction

  virtual task run();
    $display("T=%0t [Env] run task", $time);

    // Connect virtual interface handles
    d0.m_bus_vif = m_bus_vif;
    m0.m_bus_vif = m_bus_vif;

    // Connect mailboxes between each component
    d0.drv_mbx = drv_mbx;
    g0.drv_mbx = drv_mbx;

    m0.scb_mbx = scb_mbx;
    s0.scb_mbx = scb_mbx;

    // Connect event handles
    d0.drv_done = drv_done;
    g0.drv_done = drv_done;

    // Start all components - a fork join_any is used because
    // the stimulus is generated by the generator and we want the
    // simulation to exit only when the generator has finished
    // creating all transactions. Until then all other components
    // have to run in the background.

    $display("T=%0t [Env] to start fork", $time);

    fork
    	s0.run();
		  d0.run();
    	m0.run();
     	g0.run();
    join_any
  endtask
endclass
