orig/controller.sv