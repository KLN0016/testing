orig/counter.sv