orig/top_tb.sv