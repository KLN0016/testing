orig/top.sv