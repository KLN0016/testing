class fa_agt extends uvm_agent;
  `uvm_component_utils(fa_agt)

  uvm_analysis_port #(fa_tran) agt_ap;

  fa_drv drv;
  fa_mon mon;
  fa_sqr sqr;

  function new(string name, uvm_component parent);
    super.new(name, parent);
    agt_ap = new("agt_ap", this);
  endfunction

  function void build_phase(uvm_phase phase);
    super.build_phase(phase);
    mon = fa_mon::type_id::create("mon", this);
    // Only create driver and sequencer if agent is active
    if (get_is_active() == UVM_ACTIVE) begin
      drv = fa_drv::type_id::create("drv", this);
      sqr = fa_sqr::type_id::create("sqr", this);
    end
  endfunction

  function void connect_phase(uvm_phase phase);
    super.connect_phase(phase);
    // Connect monitor's analysis port to agent's analysis port
    mon.mon_ap.connect(agt_ap);
    // Connect driver to sequencer if agent active
    if (get_is_active() == UVM_ACTIVE) begin
      drv.seq_item_port.connect(sqr.seq_item_export);
    end
  endfunction
endclass
